--
-- VHDL Entity ComputerExercise1_lib.entity_name.arch_name
--
-- Created:
--          by - mfhubu.UNKNOWN (HTC219-709-SPC)
--          at - 15:25:41  4.10.2019
--
-- using Mentor Graphics HDL Designer(TM) 2019.3 (Build 4)
--
LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_arith.all;

ENTITY c1_t3_hello_led_top_level IS
   PORT( 
      btn     : IN     std_logic_vector (3 DOWNTO 0);
      sw0     : IN     std_logic;
      color   : OUT    std_logic_vector (23 DOWNTO 0);
      x_coord : OUT    std_logic_vector (7 DOWNTO 0);
      y_coord : OUT    std_logic_vector (7 DOWNTO 0)
   );

-- Declarations

END c1_t3_hello_led_top_level ;


--
-- VHDL Architecture ComputerExercise1_lib.c1_t3_hello_led_top_level.struct
--
-- Created:
--          by - mfhubu.UNKNOWN (HTC219-709-SPC)
--          at - 15:54:08  4.10.2019
--
-- Generated by Mentor Graphics' HDL Designer(TM) 2019.3 (Build 4)
--
LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_arith.all;

LIBRARY ComputerExercise1_lib;

ARCHITECTURE struct OF c1_t3_hello_led_top_level IS

   -- Architecture declarations

   -- Internal signal declarations
   SIGNAL color1    : std_logic_vector(23 DOWNTO 0);
   SIGNAL color_BGR : std_logic_vector(23 DOWNTO 0);
   SIGNAL din1      : std_logic_vector(7 DOWNTO 0);
   SIGNAL x_coord1  : std_logic_vector(7 DOWNTO 0);
   SIGNAL x_coord2  : std_logic_vector(7 DOWNTO 0);
   SIGNAL y_coord1  : std_logic_vector(7 DOWNTO 0);


   -- Component Declarations
   COMPONENT c1_t3_hello_led
   PORT (
      btn       : IN     std_logic_vector (3 DOWNTO 0);
      sw0       : IN     std_logic ;
      color_BGR : OUT    std_logic_vector (23 DOWNTO 0);
      x_coord   : OUT    std_logic_vector (7 DOWNTO 0);
      y_coord   : OUT    std_logic_vector (7 DOWNTO 0)
   );
   END COMPONENT;
   COMPONENT c1_t3_static_hello_led
   PORT (
      color   : OUT    std_logic_vector (23 DOWNTO 0);
      x_coord : OUT    std_logic_vector (7 DOWNTO 0);
      y_coord : OUT    std_logic_vector (7 DOWNTO 0)
   );
   END COMPONENT;

   -- Optional embedded configurations
   -- pragma synthesis_off
   FOR ALL : c1_t3_hello_led USE ENTITY ComputerExercise1_lib.c1_t3_hello_led;
   FOR ALL : c1_t3_static_hello_led USE ENTITY ComputerExercise1_lib.c1_t3_static_hello_led;
   -- pragma synthesis_on


BEGIN

   -- ModuleWare code(v1.12) for instance 'U_0' of 'mux'
   u_0combo_proc: PROCESS(x_coord1, x_coord2, sw0)
   BEGIN
      CASE sw0 IS
      WHEN '0' => x_coord <= x_coord1;
      WHEN '1' => x_coord <= x_coord2;
      WHEN OTHERS => x_coord <= (OTHERS => 'X');
      END CASE;
   END PROCESS u_0combo_proc;

   -- ModuleWare code(v1.12) for instance 'U_1' of 'mux'
   u_1combo_proc: PROCESS(y_coord1, din1, sw0)
   BEGIN
      CASE sw0 IS
      WHEN '0' => y_coord <= y_coord1;
      WHEN '1' => y_coord <= din1;
      WHEN OTHERS => y_coord <= (OTHERS => 'X');
      END CASE;
   END PROCESS u_1combo_proc;

   -- ModuleWare code(v1.12) for instance 'U_2' of 'mux'
   u_2combo_proc: PROCESS(color1, color_BGR, sw0)
   BEGIN
      CASE sw0 IS
      WHEN '0' => color <= color1;
      WHEN '1' => color <= color_BGR;
      WHEN OTHERS => color <= (OTHERS => 'X');
      END CASE;
   END PROCESS u_2combo_proc;

   -- Instance port mappings.
   U_3 : c1_t3_hello_led
      PORT MAP (
         btn       => btn,
         sw0       => sw0,
         color_BGR => color_BGR,
         x_coord   => x_coord2,
         y_coord   => din1
      );
   U_4 : c1_t3_static_hello_led
      PORT MAP (
         color   => color1,
         x_coord => x_coord1,
         y_coord => y_coord1
      );

END struct;
