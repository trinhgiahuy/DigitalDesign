--
-- VHDL Entity Computer_Exerccise_2_lib.C2_T3_Leftshifter.arch_name
--
-- Created:
--          by - mfhubu.UNKNOWN (HTC219-713-SPC)
--          at - 13:32:51 10.10.2019
--
-- using Mentor Graphics HDL Designer(TM) 2019.3 (Build 4)
--
LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_arith.all;

ENTITY C2_T3_Leftshifter IS
   PORT( 
      data_in  : IN     std_logic_vector (7 DOWNTO 0);
      data_out : OUT    std_logic_vector (7 DOWNTO 0)
   );

-- Declarations

END C2_T3_Leftshifter ;

