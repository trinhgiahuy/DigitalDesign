--
-- VHDL Entity Computer_Exerccise_2_lib.Half_Adder.arch_name
--
-- Created:
--          by - qkrasi.UNKNOWN (HTC219-722-SPC)
--          at - 12:09:39  8.10.2019
--
-- using Mentor Graphics HDL Designer(TM) 2019.3 (Build 4)
--
LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_arith.all;

ENTITY Half_Adder IS
   PORT( 
      x : IN     std_logic;
      y : IN     std_logic;
      c : OUT    std_logic;
      s : OUT    std_logic
   );

-- Declarations

END Half_Adder ;

