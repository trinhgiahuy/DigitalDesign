--
-- VHDL Entity ComputerExercise1_lib.entity_name.arch_name
--
-- Created:
--          by - mfhubu.UNKNOWN (HTC219-709-SPC)
--          at - 15:19:32  4.10.2019
--
-- using Mentor Graphics HDL Designer(TM) 2019.3 (Build 4)
--
LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_arith.all;

ENTITY c1_t3_static_hello_led IS
   PORT( 
      color   : OUT    std_logic_vector (23 DOWNTO 0);
      x_coord : OUT    std_logic_vector (7 DOWNTO 0);
      y_coord : OUT    std_logic_vector (7 DOWNTO 0)
   );

-- Declarations

END c1_t3_static_hello_led ;


--
-- VHDL Architecture ComputerExercise1_lib.c1_t3_static_hello_led.struct
--
-- Created:
--          by - mfhubu.UNKNOWN (HTC219-703-SPC)
--          at - 17:15:39  7.10.2019
--
-- Generated by Mentor Graphics' HDL Designer(TM) 2019.3 (Build 4)
--
LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_arith.all;


ARCHITECTURE struct OF c1_t3_static_hello_led IS

   -- Architecture declarations

   -- Internal signal declarations



BEGIN

   -- ModuleWare code(v1.12) for instance 'U_0' of 'constval'
   x_coord <= "00100000";

   -- ModuleWare code(v1.12) for instance 'U_1' of 'constval'
   y_coord <= "00100000";

   -- ModuleWare code(v1.12) for instance 'U_2' of 'constval'
   color <= "000000000000010010110000";

   -- Instance port mappings.

END struct;
