--* ><(((('> * Puli puli * ><(((('> // Ƹ̵̡Ӝ̵̨̄Ʒ * swish swish* Ƹ̵̡Ӝ̵̨̄Ʒ Ƹ̵̡Ӝ̵̨̄Ʒ // (っ◕‿◕)╭∩╮^H^H^Hっ
LIBRARY ieee;USE ieee.std_logic_1164.all;USE ieee.std_logic_arith.all;ENTITY reg_bank_64px IS PORT(clk:IN std_logic;nullify:IN std_logic;zd58ce0c39:IN std_logic_vector(23 DOWNTO 0);rst_n:IN std_logic;write:IN std_logic;x:IN std_logic_vector(7 DOWNTO 0);y:IN std_logic_vector(7 DOWNTO 0);pix_out:OUT std_logic_vector(23 DOWNTO 0));END reg_bank_64px ;LIBRARY ieee;USE ieee.std_logic_1164.all;USE ieee.std_logic_arith.all;LIBRARY Computer_Exercise_5_lib;ARCHITECTURE struct OF reg_bank_64px IS SIGNAL z508ec0017:std_logic;SIGNAL z1934d98a3:std_logic;SIGNAL zb48298c48:std_logic;SIGNAL z9f041aaff:std_logic;SIGNAL zcf058ee7c:std_logic;SIGNAL ze6d31b4ac:std_logic;SIGNAL z1b791bfd5:std_logic;SIGNAL z45a1dff88:std_logic;SIGNAL zc83e54d35:std_logic_vector(2 DOWNTO 0);SIGNAL z22f92b4dd:std_logic;SIGNAL z75dc1577a:std_logic;SIGNAL z833ab3bd5:std_logic;SIGNAL zc57c46db4:std_logic;SIGNAL z1ea89dc0d:std_logic;SIGNAL zcd48e1f4f:std_logic;SIGNAL z36424fa31:std_logic;SIGNAL z0068e7d64:std_logic;SIGNAL zb30429bb4:std_logic;SIGNAL z36f79a239:std_logic_vector(3 DOWNTO 0);SIGNAL pixd_out:std_logic_vector(23 DOWNTO 0);SIGNAL z564ee05a3:std_logic_vector(23 DOWNTO 0);SIGNAL z0a9315da3:std_logic_vector(23 DOWNTO 0);SIGNAL z6bb6c7052:std_logic_vector(23 DOWNTO 0);SIGNAL z163c5325c:std_logic_vector(23 DOWNTO 0);SIGNAL z84b2eb77e:std_logic_vector(23 DOWNTO 0);SIGNAL zed22165f2:std_logic_vector(23 DOWNTO 0);SIGNAL z90a7dbf30:std_logic_vector(23 DOWNTO 0);SIGNAL zf090fac59:std_logic_vector(7 DOWNTO 0);COMPONENT reg_bank_1col PORT(clk:IN std_logic ;nullify:IN std_logic ;pixd_in:IN std_logic_vector(23 DOWNTO 0);rst_n:IN std_logic ;write:IN std_logic ;y:IN std_logic_vector(7 DOWNTO 0);pixd_out:OUT std_logic_vector(23 DOWNTO 0));END COMPONENT;FOR ALL:reg_bank_1col USE ENTITY Computer_Exercise_5_lib.reg_bank_1col;BEGIN z508ec0017<=write AND z1934d98a3;zb48298c48<=write AND z0068e7d64;z75dc1577a<=write AND zb30429bb4;z833ab3bd5<=write AND z9f041aaff;zc57c46db4<=write AND zcf058ee7c;z1ea89dc0d<=write AND ze6d31b4ac;zcd48e1f4f<=write AND z1b791bfd5;z36424fa31<=write AND z45a1dff88;z22f92b4dd<='1';zd4351336a:PROCESS(z22f92b4dd, x)BEGIN IF(x(0)=z22f92b4dd)THEN z36f79a239<="0000";ELSIF(x(1)=z22f92b4dd)THEN z36f79a239<="0001";ELSIF(x(2)=z22f92b4dd)THEN z36f79a239<="0010";ELSIF(x(3)=z22f92b4dd)THEN z36f79a239<="0011";ELSIF(x(4)=z22f92b4dd)THEN z36f79a239<="0100";ELSIF(x(5)=z22f92b4dd)THEN z36f79a239<="0101";ELSIF(x(6)=z22f92b4dd)THEN z36f79a239<="0110";ELSIF(x(7)=z22f92b4dd)THEN z36f79a239<="0111";ELSE z36f79a239<="1000";END IF;END PROCESS zd4351336a;zc83e54d35<=z36f79a239(2)& z36f79a239(1)& z36f79a239(0);z16921971f:PROCESS(pixd_out, z564ee05a3, z0a9315da3, z6bb6c7052, z163c5325c, z84b2eb77e, zed22165f2, z90a7dbf30, zc83e54d35)BEGIN CASE zc83e54d35 IS WHEN"000"=>pix_out<=pixd_out;WHEN"001"=>pix_out<=z564ee05a3;WHEN"010"=>pix_out<=z0a9315da3;WHEN"011"=>pix_out<=z6bb6c7052;WHEN"100"=>pix_out<=z163c5325c;WHEN"101"=>pix_out<=z84b2eb77e;WHEN"110"=>pix_out<=zed22165f2;WHEN"111"=>pix_out<=z90a7dbf30;WHEN OTHERS=>pix_out<=(OTHERS=>'X');END CASE;END PROCESS z16921971f;zf090fac59<=x;z193f2f0f4:PROCESS(zf090fac59)VARIABLE z925f2bf10:std_logic_vector(7 DOWNTO 0);BEGIN z925f2bf10:=zf090fac59(7 DOWNTO 0);z1934d98a3<=z925f2bf10(0);z0068e7d64<=z925f2bf10(1);zb30429bb4<=z925f2bf10(2);z9f041aaff<=z925f2bf10(3);zcf058ee7c<=z925f2bf10(4);ze6d31b4ac<=z925f2bf10(5);z1b791bfd5<=z925f2bf10(6);z45a1dff88<=z925f2bf10(7);END PROCESS z193f2f0f4;U_0:reg_bank_1col PORT MAP(clk=>clk,nullify=>nullify,pixd_in=>zd58ce0c39,rst_n=>rst_n,write=>z508ec0017,y=>y,pixd_out=>pixd_out);U_1:reg_bank_1col PORT MAP(clk=>clk,nullify=>nullify,pixd_in=>zd58ce0c39,rst_n=>rst_n,write=>zb48298c48,y=>y,pixd_out=>z564ee05a3);U_2:reg_bank_1col PORT MAP(clk=>clk,nullify=>nullify,pixd_in=>zd58ce0c39,rst_n=>rst_n,write=>z75dc1577a,y=>y,pixd_out=>z0a9315da3);U_3:reg_bank_1col PORT MAP(clk=>clk,nullify=>nullify,pixd_in=>zd58ce0c39,rst_n=>rst_n,write=>z833ab3bd5,y=>y,pixd_out=>z6bb6c7052);U_4:reg_bank_1col PORT MAP(clk=>clk,nullify=>nullify,pixd_in=>zd58ce0c39,rst_n=>rst_n,write=>zc57c46db4,y=>y,pixd_out=>z163c5325c);U_5:reg_bank_1col PORT MAP(clk=>clk,nullify=>nullify,pixd_in=>zd58ce0c39,rst_n=>rst_n,write=>z1ea89dc0d,y=>y,pixd_out=>z84b2eb77e);U_6:reg_bank_1col PORT MAP(clk=>clk,nullify=>nullify,pixd_in=>zd58ce0c39,rst_n=>rst_n,write=>zcd48e1f4f,y=>y,pixd_out=>zed22165f2);U_7:reg_bank_1col PORT MAP(clk=>clk,nullify=>nullify,pixd_in=>zd58ce0c39,rst_n=>rst_n,write=>z36424fa31,y=>y,pixd_out=>z90a7dbf30);END struct;