--
-- VHDL Entity Computer_Exerccise_2_lib.C2_T2_Decrementer.arch_name
--
-- Created:
--          by - qkrasi.UNKNOWN (HTC219-722-SPC)
--          at - 12:54:59  8.10.2019
--
-- using Mentor Graphics HDL Designer(TM) 2019.3 (Build 4)
--
LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_arith.all;

ENTITY C2_T2_Decrementer IS
   PORT( 
      Input  : IN     std_logic_vector (2 DOWNTO 0);
      Output : OUT    std_logic_vector (2 DOWNTO 0)
   );

-- Declarations

END C2_T2_Decrementer ;

