--
-- VHDL Entity Computer_Exerccise_2_lib.C2_T7_Basic_Alien.arch_name
--
-- Created:
--          by - mfhubu.UNKNOWN (HTC219-711-SPC)
--          at - 11:22:06 11.10.2019
--
-- using Mentor Graphics HDL Designer(TM) 2019.3 (Build 4)
--
LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_arith.all;

ENTITY C2_T7_Basic_Alien IS
   PORT( 
      clk         : IN     std_logic;
      enable      : IN     std_logic;
      enable_slow : IN     std_logic;
      hit         : IN     std_logic;
      rst_n       : IN     std_logic;
      speed       : IN     std_logic;
      alien_col   : OUT    std_logic_vector (23 DOWNTO 0);
      x_coord     : OUT    std_logic_vector (7 DOWNTO 0);
      y_coord     : OUT    std_logic_vector (7 DOWNTO 0)
   );

-- Declarations

END C2_T7_Basic_Alien ;


--
-- VHDL Architecture Computer_Exerccise_2_lib.C2_T7_Basic_Alien.struct
--
-- Created:
--          by - mfhubu.UNKNOWN (HTC219-708-SPC)
--          at - 11:43:43 19.11.2019
--
-- Generated by Mentor Graphics' HDL Designer(TM) 2019.3 (Build 4)
--
LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_arith.all;

LIBRARY Computer_Exerccise_2_lib;

ARCHITECTURE struct OF C2_T7_Basic_Alien IS

   -- Architecture declarations

   -- Internal signal declarations
   SIGNAL data_out : std_logic_vector(7 DOWNTO 0);
   SIGNAL din2     : std_logic_vector(7 DOWNTO 0);
   SIGNAL dout3    : std_logic_vector(7 DOWNTO 0);
   SIGNAL dout6    : std_logic_vector(1 DOWNTO 0);
   SIGNAL enable1  : std_logic;

   -- Implicit buffer signal declarations
   SIGNAL x_coord_internal : std_logic_vector (7 DOWNTO 0);


   -- ModuleWare signal declarations(v1.12) for instance 'U_1' of 'adff'
   SIGNAL mw_U_1reg_cval : std_logic_vector(7 DOWNTO 0);

   -- Component Declarations
   COMPONENT Basic_Alien_Direction
   PORT (
      clk       : IN     std_logic ;
      enable    : IN     std_logic ;
      rst_n     : IN     std_logic ;
      x_0       : IN     std_logic ;                   -- Condition TO switch direction
      x_7       : IN     std_logic ;                   -- Condition TO switch direction
      direction : OUT    std_logic_vector (1 DOWNTO 0) -- 2 MSB allow TO shift - 2 LSB decide direction
   );
   END COMPONENT;
   COMPONENT Basic_Alien_color
   PORT (
      clk       : IN     std_logic ;
      hit       : IN     std_logic ;
      rst_n     : IN     std_logic ;
      alien_col : OUT    std_logic_vector (23 DOWNTO 0)
   );
   END COMPONENT;
   COMPONENT Basic_Alien_y_coord
   PORT (
      clk     : IN     std_logic ;
      rst_n   : IN     std_logic ;
      y_coord : OUT    std_logic_vector (7 DOWNTO 0)
   );
   END COMPONENT;
   COMPONENT C2_T3_Leftshifter
   PORT (
      data_in  : IN     std_logic_vector (7 DOWNTO 0);
      data_out : OUT    std_logic_vector (7 DOWNTO 0)
   );
   END COMPONENT;
   COMPONENT C2_T4_Rightshifter
   PORT (
      x : IN     std_logic_vector (7 DOWNTO 0);
      y : OUT    std_logic_vector (7 DOWNTO 0)
   );
   END COMPONENT;

   -- Optional embedded configurations
   -- pragma synthesis_off
   FOR ALL : Basic_Alien_Direction USE ENTITY Computer_Exerccise_2_lib.Basic_Alien_Direction;
   FOR ALL : Basic_Alien_color USE ENTITY Computer_Exerccise_2_lib.Basic_Alien_color;
   FOR ALL : Basic_Alien_y_coord USE ENTITY Computer_Exerccise_2_lib.Basic_Alien_y_coord;
   FOR ALL : C2_T3_Leftshifter USE ENTITY Computer_Exerccise_2_lib.C2_T3_Leftshifter;
   FOR ALL : C2_T4_Rightshifter USE ENTITY Computer_Exerccise_2_lib.C2_T4_Rightshifter;
   -- pragma synthesis_on


BEGIN

   -- ModuleWare code(v1.12) for instance 'U_1' of 'adff'
   x_coord_internal <= mw_U_1reg_cval;
   u_1seq_proc: PROCESS (clk, rst_n)
   BEGIN
      IF (rst_n = '0') THEN
         mw_U_1reg_cval <= "00100000";
      ELSIF (clk'EVENT AND clk='1') THEN
         mw_U_1reg_cval <= dout3;
      END IF;
   END PROCESS u_1seq_proc;

   -- ModuleWare code(v1.12) for instance 'U_3' of 'mux'
   u_3combo_proc: PROCESS(enable_slow, enable, speed)
   BEGIN
      CASE speed IS
      WHEN '0' => enable1 <= enable_slow;
      WHEN '1' => enable1 <= enable;
      WHEN OTHERS => enable1 <= 'X';
      END CASE;
   END PROCESS u_3combo_proc;

   -- ModuleWare code(v1.12) for instance 'U_16' of 'mux'
   u_16combo_proc: PROCESS(x_coord_internal, data_out, din2, dout6)
   BEGIN
      CASE dout6 IS
      WHEN "00" => dout3 <= x_coord_internal;
      WHEN "01" => dout3 <= data_out;
      WHEN "10" => dout3 <= din2;
      WHEN "11" => dout3 <= x_coord_internal;
      WHEN OTHERS => dout3 <= (OTHERS => 'X');
      END CASE;
   END PROCESS u_16combo_proc;

   -- Instance port mappings.
   U_2 : Basic_Alien_Direction
      PORT MAP (
         clk       => clk,
         enable    => enable1,
         rst_n     => rst_n,
         x_0       => x_coord_internal(0),
         x_7       => x_coord_internal(7),
         direction => dout6
      );
   U_0 : Basic_Alien_color
      PORT MAP (
         clk       => clk,
         hit       => hit,
         rst_n     => rst_n,
         alien_col => alien_col
      );
   U_4 : Basic_Alien_y_coord
      PORT MAP (
         clk     => clk,
         rst_n   => rst_n,
         y_coord => y_coord
      );
   U_8 : C2_T3_Leftshifter
      PORT MAP (
         data_in  => x_coord_internal,
         data_out => data_out
      );
   U_7 : C2_T4_Rightshifter
      PORT MAP (
         x => x_coord_internal,
         y => din2
      );

   -- Implicit buffered output assignments
   x_coord <= x_coord_internal;

END struct;
